`default_nettype none

// Utility module aliases for IP compatibility

module ef_util_ned (
    input wire clk,
    input wire in,
    output wire out
);
    aucohl_ned ned_inst (.clk(clk), .in(in), .out(out));
endmodule

module cf_util_ped (
    input wire clk,
    input wire in,
    output wire out
);
    aucohl_ped ped_inst (.clk(clk), .in(in), .out(out));
endmodule

module cf_util_fifo #(parameter DW = 8, AW = 4) (
    input wire clk,
    input wire rst_n,
    input wire rd,
    input wire wr,
    input wire flush,
    input wire [DW-1:0] wdata,
    output wire empty,
    output wire full,
    output wire [DW-1:0] rdata,
    output wire [AW-1:0] level
);
    aucohl_fifo #(.DW(DW), .AW(AW)) fifo_inst (
        .clk(clk),
        .rst_n(rst_n),
        .rd(rd),
        .wr(wr),
        .flush(flush),
        .wdata(wdata),
        .empty(empty),
        .full(full),
        .rdata(rdata),
        .level(level)
    );
endmodule

module ef_util_gating_cell (
    input wire clk,
    input wire clk_en,
    output wire clk_o
);
    ef_gating_cell gating_inst (
        .clk(clk), 
        .rst_n(1'b1), 
        .clk_en(clk_en), 
        .clk_o(clk_o)
    );
endmodule

module cf_util_gating_cell (
    input wire clk,
    input wire clk_en,
    output wire clk_o
);
    ef_gating_cell gating_inst (
        .clk(clk), 
        .rst_n(1'b1), 
        .clk_en(clk_en), 
        .clk_o(clk_o)
    );
endmodule

module ef_util_sync #(parameter NUM_STAGES = 2) (
    input wire clk,
    input wire in,
    output wire out
);
    aucohl_sync #(.NUM_STAGES(NUM_STAGES)) sync_inst (.clk(clk), .in(in), .out(out));
endmodule

module ef_util_ped (
    input wire clk,
    input wire in,
    output wire out
);
    aucohl_ped ped_inst (.clk(clk), .in(in), .out(out));
endmodule

`default_nettype wire